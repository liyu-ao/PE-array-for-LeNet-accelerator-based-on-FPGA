module add(
    input  [15:0] A,
    input  [15:0] B,
    output  [15:0] out
);
    wire [15:0] x,y,sum;

    assign x=(A[15]==1)?(((A[14:0])==15'b0)?{16'b00000000}:{1'b1,~A[14:0]+1'b1}):({A[15:0]});
    assign y=(B[15]==1)?(((B[14:0])==15'b0)?{16'b00000000}:{1'b1,~B[14:0]+1'b1}):({B[15:0]});//当输入是10000000时转换为00000000参与计算

    assign sum = x + y;

    assign out = (x[15] & y[15])?  {1'b1,~sum[14:0]+1'b1}: //两个负数
                    ( (x[15] || y[15])?(sum[15]?{1'b1,~sum[14:0]+1'b1}:{1'b0,sum[14:0]}): //一正一负 
						{1'b0,sum[14:0]} );	// （两个正数）  	

endmodule 
